/*************************************************************************
 > Copyright (C) 2021 Sangfor Ltd. All rights reserved.
 > File Name   : defines.sv
 > Author      : bhyou
 > Mail        : bhyou@foxmail.com 
 > Created Time: Wed 07 Jul 2021 07:52:07 PM CST
 ************************************************************************/

 
`define DEBUG_MEDIUM
`define CollectRadius 25
`define LocalThreshold 5
`define SummingThreshold 15
 
 //`define testingDiscriminator
//`define testingAnalogFrontend
// `define testingPixelCells
// `define testingPixelArray
// `define testingChannel
//`define testAnalogFrontEnd
//`define testingAnalogFrontendArray
 `define testAnalogEnvironment